library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity Test_CDC2 is
end Test_CDC2;

architecture Behavioral of Test_CDC2 is
    component Main
        Port (
              -- Switch
              e1 : in STD_LOGIC;
              e2 : in STD_LOGIC;
              e11 : in STD_LOGIC; -- And
              e12 : in STD_LOGIC; -- Or
              e13 : in STD_LOGIC; -- Not
              e14 : in STD_LOGIC; -- Xor
              e15 : in STD_LOGIC; -- Nand
              e16 : in STD_LOGIC; -- Nor
              
              -- LED
              l1 : out STD_LOGIC;
              l2 : out STD_LOGIC;
              l11 : out STD_LOGIC;
              l12 : out STD_LOGIC;
              l13 : out STD_LOGIC;
              l14 : out STD_LOGIC;
              l15 : out STD_LOGIC;
              l16 : out STD_LOGIC;
              
              -- Display Bloc
              a : out STD_LOGIC;
              b : out STD_LOGIC;
              c : out STD_LOGIC;
              d : out STD_LOGIC;
              e : out STD_LOGIC;
              f : out STD_LOGIC;
              g : out STD_LOGIC;
              dp : out STD_LOGIC);
    end component;
    
    signal e1: STD_LOGIC:='0';
    signal e2: STD_LOGIC:='0';
    signal e11: STD_LOGIC:='0';
    signal e12: STD_LOGIC:='0';
    signal e13: STD_LOGIC:='0';
    signal e14: STD_LOGIC:='0';
    signal e15: STD_LOGIC:='0';
    signal e16: STD_LOGIC:='0';
    signal l1: STD_LOGIC:='0';
    signal l2: STD_LOGIC:='0';
    signal l11: STD_LOGIC:='0';
    signal l12: STD_LOGIC:='0';
    signal l13: STD_LOGIC:='0';
    signal l14: STD_LOGIC:='0';
    signal l15: STD_LOGIC:='0';
    signal l16: STD_LOGIC:='0';
    signal a: STD_LOGIC;
    signal b: STD_LOGIC;
    signal c: STD_LOGIC;
    signal d: STD_LOGIC;
    signal e: STD_LOGIC;
    signal f: STD_LOGIC;
    signal g: STD_LOGIC;
    signal dp : STD_Logic;
    
    constant period:time :=2 ns;
begin
    Generate_In: process
            begin
            e11 <='0'; e12 <='0'; e13 <='0'; e14 <='0'; e15 <='0'; e16 <='0'; e1 <='0'; e2 <='0'; wait for period;
            e11 <='1'; e12 <='0'; e13 <='0'; e14 <='0'; e15 <='0'; e16 <='0'; e1 <='0'; e2 <='0'; wait for period;
            e11 <='0'; e12 <='1'; e13 <='0'; e14 <='0'; e15 <='0'; e16 <='0'; e1 <='0'; e2 <='0'; wait for period;
            e11 <='1'; e12 <='1'; e13 <='0'; e14 <='0'; e15 <='0'; e16 <='0'; e1 <='0'; e2 <='0'; wait for period;
            e11 <='0'; e12 <='0'; e13 <='1'; e14 <='0'; e15 <='0'; e16 <='0'; e1 <='0'; e2 <='0'; wait for period;
            e11 <='1'; e12 <='0'; e13 <='1'; e14 <='0'; e15 <='0'; e16 <='0'; e1 <='0'; e2 <='0'; wait for period;
            e11 <='0'; e12 <='1'; e13 <='1'; e14 <='0'; e15 <='0'; e16 <='0'; e1 <='0'; e2 <='0'; wait for period;
            e11 <='1'; e12 <='1'; e13 <='1'; e14 <='0'; e15 <='0'; e16 <='0'; e1 <='0'; e2 <='0'; wait for period;
            e11 <='0'; e12 <='0'; e13 <='0'; e14 <='1'; e15 <='0'; e16 <='0'; e1 <='0'; e2 <='0'; wait for period;
            e11 <='1'; e12 <='0'; e13 <='0'; e14 <='1'; e15 <='0'; e16 <='0'; e1 <='0'; e2 <='0'; wait for period;
            e11 <='0'; e12 <='1'; e13 <='0'; e14 <='1'; e15 <='0'; e16 <='0'; e1 <='0'; e2 <='0'; wait for period;
            e11 <='1'; e12 <='1'; e13 <='0'; e14 <='1'; e15 <='0'; e16 <='0'; e1 <='0'; e2 <='0'; wait for period;
            e11 <='0'; e12 <='0'; e13 <='1'; e14 <='1'; e15 <='0'; e16 <='0'; e1 <='0'; e2 <='0'; wait for period;
            e11 <='1'; e12 <='0'; e13 <='1'; e14 <='1'; e15 <='0'; e16 <='0'; e1 <='0'; e2 <='0'; wait for period;
            e11 <='0'; e12 <='1'; e13 <='1'; e14 <='1'; e15 <='0'; e16 <='0'; e1 <='0'; e2 <='0'; wait for period;
            e11 <='1'; e12 <='1'; e13 <='1'; e14 <='1'; e15 <='0'; e16 <='0'; e1 <='0'; e2 <='0'; wait for period;
            e11 <='0'; e12 <='0'; e13 <='0'; e14 <='0'; e15 <='1'; e16 <='0'; e1 <='0'; e2 <='0'; wait for period;
            e11 <='1'; e12 <='0'; e13 <='0'; e14 <='0'; e15 <='1'; e16 <='0'; e1 <='0'; e2 <='0'; wait for period;
            e11 <='0'; e12 <='1'; e13 <='0'; e14 <='0'; e15 <='1'; e16 <='0'; e1 <='0'; e2 <='0'; wait for period;
            e11 <='1'; e12 <='1'; e13 <='0'; e14 <='0'; e15 <='1'; e16 <='0'; e1 <='0'; e2 <='0'; wait for period;
            e11 <='0'; e12 <='0'; e13 <='1'; e14 <='0'; e15 <='1'; e16 <='0'; e1 <='0'; e2 <='0'; wait for period;
            e11 <='1'; e12 <='0'; e13 <='1'; e14 <='0'; e15 <='1'; e16 <='0'; e1 <='0'; e2 <='0'; wait for period;
            e11 <='0'; e12 <='1'; e13 <='1'; e14 <='0'; e15 <='1'; e16 <='0'; e1 <='0'; e2 <='0'; wait for period;
            e11 <='1'; e12 <='1'; e13 <='1'; e14 <='0'; e15 <='1'; e16 <='0'; e1 <='0'; e2 <='0'; wait for period;
            e11 <='0'; e12 <='0'; e13 <='0'; e14 <='1'; e15 <='1'; e16 <='0'; e1 <='0'; e2 <='0'; wait for period;
            e11 <='1'; e12 <='0'; e13 <='0'; e14 <='1'; e15 <='1'; e16 <='0'; e1 <='0'; e2 <='0'; wait for period;
            e11 <='0'; e12 <='1'; e13 <='0'; e14 <='1'; e15 <='1'; e16 <='0'; e1 <='0'; e2 <='0'; wait for period;
            e11 <='1'; e12 <='1'; e13 <='0'; e14 <='1'; e15 <='1'; e16 <='0'; e1 <='0'; e2 <='0'; wait for period;
            e11 <='0'; e12 <='0'; e13 <='1'; e14 <='1'; e15 <='1'; e16 <='0'; e1 <='0'; e2 <='0'; wait for period;
            e11 <='1'; e12 <='0'; e13 <='1'; e14 <='1'; e15 <='1'; e16 <='0'; e1 <='0'; e2 <='0'; wait for period;
            e11 <='0'; e12 <='1'; e13 <='1'; e14 <='1'; e15 <='1'; e16 <='0'; e1 <='0'; e2 <='0'; wait for period;
            e11 <='1'; e12 <='1'; e13 <='1'; e14 <='1'; e15 <='1'; e16 <='0'; e1 <='0'; e2 <='0'; wait for period;
            e11 <='0'; e12 <='0'; e13 <='0'; e14 <='0'; e15 <='0'; e16 <='1'; e1 <='0'; e2 <='0'; wait for period;
            e11 <='1'; e12 <='0'; e13 <='0'; e14 <='0'; e15 <='0'; e16 <='1'; e1 <='0'; e2 <='0'; wait for period;
            e11 <='0'; e12 <='1'; e13 <='0'; e14 <='0'; e15 <='0'; e16 <='1'; e1 <='0'; e2 <='0'; wait for period;
            e11 <='1'; e12 <='1'; e13 <='0'; e14 <='0'; e15 <='0'; e16 <='1'; e1 <='0'; e2 <='0'; wait for period;
            e11 <='0'; e12 <='0'; e13 <='1'; e14 <='0'; e15 <='0'; e16 <='1'; e1 <='0'; e2 <='0'; wait for period;
            e11 <='1'; e12 <='0'; e13 <='1'; e14 <='0'; e15 <='0'; e16 <='1'; e1 <='0'; e2 <='0'; wait for period;
            e11 <='0'; e12 <='1'; e13 <='1'; e14 <='0'; e15 <='0'; e16 <='1'; e1 <='0'; e2 <='0'; wait for period;
            e11 <='1'; e12 <='1'; e13 <='1'; e14 <='0'; e15 <='0'; e16 <='1'; e1 <='0'; e2 <='0'; wait for period;
            e11 <='0'; e12 <='0'; e13 <='0'; e14 <='1'; e15 <='0'; e16 <='1'; e1 <='0'; e2 <='0'; wait for period;
            e11 <='1'; e12 <='0'; e13 <='0'; e14 <='1'; e15 <='0'; e16 <='1'; e1 <='0'; e2 <='0'; wait for period;
            e11 <='0'; e12 <='1'; e13 <='0'; e14 <='1'; e15 <='0'; e16 <='1'; e1 <='0'; e2 <='0'; wait for period;
            e11 <='1'; e12 <='1'; e13 <='0'; e14 <='1'; e15 <='0'; e16 <='1'; e1 <='0'; e2 <='0'; wait for period;
            e11 <='0'; e12 <='0'; e13 <='1'; e14 <='1'; e15 <='0'; e16 <='1'; e1 <='0'; e2 <='0'; wait for period;
            e11 <='1'; e12 <='0'; e13 <='1'; e14 <='1'; e15 <='0'; e16 <='1'; e1 <='0'; e2 <='0'; wait for period;
            e11 <='0'; e12 <='1'; e13 <='1'; e14 <='1'; e15 <='0'; e16 <='1'; e1 <='0'; e2 <='0'; wait for period;
            e11 <='1'; e12 <='1'; e13 <='1'; e14 <='1'; e15 <='0'; e16 <='1'; e1 <='0'; e2 <='0'; wait for period;
            e11 <='0'; e12 <='0'; e13 <='0'; e14 <='0'; e15 <='1'; e16 <='1'; e1 <='0'; e2 <='0'; wait for period;
            e11 <='1'; e12 <='0'; e13 <='0'; e14 <='0'; e15 <='1'; e16 <='1'; e1 <='0'; e2 <='0'; wait for period;
            e11 <='0'; e12 <='1'; e13 <='0'; e14 <='0'; e15 <='1'; e16 <='1'; e1 <='0'; e2 <='0'; wait for period;
            e11 <='1'; e12 <='1'; e13 <='0'; e14 <='0'; e15 <='1'; e16 <='1'; e1 <='0'; e2 <='0'; wait for period;
            e11 <='0'; e12 <='0'; e13 <='1'; e14 <='0'; e15 <='1'; e16 <='1'; e1 <='0'; e2 <='0'; wait for period;
            e11 <='1'; e12 <='0'; e13 <='1'; e14 <='0'; e15 <='1'; e16 <='1'; e1 <='0'; e2 <='0'; wait for period;
            e11 <='0'; e12 <='1'; e13 <='1'; e14 <='0'; e15 <='1'; e16 <='1'; e1 <='0'; e2 <='0'; wait for period;
            e11 <='1'; e12 <='1'; e13 <='1'; e14 <='0'; e15 <='1'; e16 <='1'; e1 <='0'; e2 <='0'; wait for period;
            e11 <='0'; e12 <='0'; e13 <='0'; e14 <='1'; e15 <='1'; e16 <='1'; e1 <='0'; e2 <='0'; wait for period;
            e11 <='1'; e12 <='0'; e13 <='0'; e14 <='1'; e15 <='1'; e16 <='1'; e1 <='0'; e2 <='0'; wait for period;
            e11 <='0'; e12 <='1'; e13 <='0'; e14 <='1'; e15 <='1'; e16 <='1'; e1 <='0'; e2 <='0'; wait for period;
            e11 <='1'; e12 <='1'; e13 <='0'; e14 <='1'; e15 <='1'; e16 <='1'; e1 <='0'; e2 <='0'; wait for period;
            e11 <='0'; e12 <='0'; e13 <='1'; e14 <='1'; e15 <='1'; e16 <='1'; e1 <='0'; e2 <='0'; wait for period;
            e11 <='1'; e12 <='0'; e13 <='1'; e14 <='1'; e15 <='1'; e16 <='1'; e1 <='0'; e2 <='0'; wait for period;
            e11 <='0'; e12 <='1'; e13 <='1'; e14 <='1'; e15 <='1'; e16 <='1'; e1 <='0'; e2 <='0'; wait for period;
            e11 <='1'; e12 <='1'; e13 <='1'; e14 <='1'; e15 <='1'; e16 <='1'; e1 <='0'; e2 <='0'; wait for period;
            e11 <='0'; e12 <='0'; e13 <='0'; e14 <='0'; e15 <='0'; e16 <='0'; e1 <='1'; e2 <='0'; wait for period;
            e11 <='1'; e12 <='0'; e13 <='0'; e14 <='0'; e15 <='0'; e16 <='0'; e1 <='1'; e2 <='0'; wait for period;
            e11 <='0'; e12 <='1'; e13 <='0'; e14 <='0'; e15 <='0'; e16 <='0'; e1 <='1'; e2 <='0'; wait for period;
            e11 <='1'; e12 <='1'; e13 <='0'; e14 <='0'; e15 <='0'; e16 <='0'; e1 <='1'; e2 <='0'; wait for period;
            e11 <='0'; e12 <='0'; e13 <='1'; e14 <='0'; e15 <='0'; e16 <='0'; e1 <='1'; e2 <='0'; wait for period;
            e11 <='1'; e12 <='0'; e13 <='1'; e14 <='0'; e15 <='0'; e16 <='0'; e1 <='1'; e2 <='0'; wait for period;
            e11 <='0'; e12 <='1'; e13 <='1'; e14 <='0'; e15 <='0'; e16 <='0'; e1 <='1'; e2 <='0'; wait for period;
            e11 <='1'; e12 <='1'; e13 <='1'; e14 <='0'; e15 <='0'; e16 <='0'; e1 <='1'; e2 <='0'; wait for period;
            e11 <='0'; e12 <='0'; e13 <='0'; e14 <='1'; e15 <='0'; e16 <='0'; e1 <='1'; e2 <='0'; wait for period;
            e11 <='1'; e12 <='0'; e13 <='0'; e14 <='1'; e15 <='0'; e16 <='0'; e1 <='1'; e2 <='0'; wait for period;
            e11 <='0'; e12 <='1'; e13 <='0'; e14 <='1'; e15 <='0'; e16 <='0'; e1 <='1'; e2 <='0'; wait for period;
            e11 <='1'; e12 <='1'; e13 <='0'; e14 <='1'; e15 <='0'; e16 <='0'; e1 <='1'; e2 <='0'; wait for period;
            e11 <='0'; e12 <='0'; e13 <='1'; e14 <='1'; e15 <='0'; e16 <='0'; e1 <='1'; e2 <='0'; wait for period;
            e11 <='1'; e12 <='0'; e13 <='1'; e14 <='1'; e15 <='0'; e16 <='0'; e1 <='1'; e2 <='0'; wait for period;
            e11 <='0'; e12 <='1'; e13 <='1'; e14 <='1'; e15 <='0'; e16 <='0'; e1 <='1'; e2 <='0'; wait for period;
            e11 <='1'; e12 <='1'; e13 <='1'; e14 <='1'; e15 <='0'; e16 <='0'; e1 <='1'; e2 <='0'; wait for period;
            e11 <='0'; e12 <='0'; e13 <='0'; e14 <='0'; e15 <='1'; e16 <='0'; e1 <='1'; e2 <='0'; wait for period;
            e11 <='1'; e12 <='0'; e13 <='0'; e14 <='0'; e15 <='1'; e16 <='0'; e1 <='1'; e2 <='0'; wait for period;
            e11 <='0'; e12 <='1'; e13 <='0'; e14 <='0'; e15 <='1'; e16 <='0'; e1 <='1'; e2 <='0'; wait for period;
            e11 <='1'; e12 <='1'; e13 <='0'; e14 <='0'; e15 <='1'; e16 <='0'; e1 <='1'; e2 <='0'; wait for period;
            e11 <='0'; e12 <='0'; e13 <='1'; e14 <='0'; e15 <='1'; e16 <='0'; e1 <='1'; e2 <='0'; wait for period;
            e11 <='1'; e12 <='0'; e13 <='1'; e14 <='0'; e15 <='1'; e16 <='0'; e1 <='1'; e2 <='0'; wait for period;
            e11 <='0'; e12 <='1'; e13 <='1'; e14 <='0'; e15 <='1'; e16 <='0'; e1 <='1'; e2 <='0'; wait for period;
            e11 <='1'; e12 <='1'; e13 <='1'; e14 <='0'; e15 <='1'; e16 <='0'; e1 <='1'; e2 <='0'; wait for period;
            e11 <='0'; e12 <='0'; e13 <='0'; e14 <='1'; e15 <='1'; e16 <='0'; e1 <='1'; e2 <='0'; wait for period;
            e11 <='1'; e12 <='0'; e13 <='0'; e14 <='1'; e15 <='1'; e16 <='0'; e1 <='1'; e2 <='0'; wait for period;
            e11 <='0'; e12 <='1'; e13 <='0'; e14 <='1'; e15 <='1'; e16 <='0'; e1 <='1'; e2 <='0'; wait for period;
            e11 <='1'; e12 <='1'; e13 <='0'; e14 <='1'; e15 <='1'; e16 <='0'; e1 <='1'; e2 <='0'; wait for period;
            e11 <='0'; e12 <='0'; e13 <='1'; e14 <='1'; e15 <='1'; e16 <='0'; e1 <='1'; e2 <='0'; wait for period;
            e11 <='1'; e12 <='0'; e13 <='1'; e14 <='1'; e15 <='1'; e16 <='0'; e1 <='1'; e2 <='0'; wait for period;
            e11 <='0'; e12 <='1'; e13 <='1'; e14 <='1'; e15 <='1'; e16 <='0'; e1 <='1'; e2 <='0'; wait for period;
            e11 <='1'; e12 <='1'; e13 <='1'; e14 <='1'; e15 <='1'; e16 <='0'; e1 <='1'; e2 <='0'; wait for period;
            e11 <='0'; e12 <='0'; e13 <='0'; e14 <='0'; e15 <='0'; e16 <='1'; e1 <='1'; e2 <='0'; wait for period;
            e11 <='1'; e12 <='0'; e13 <='0'; e14 <='0'; e15 <='0'; e16 <='1'; e1 <='1'; e2 <='0'; wait for period;
            e11 <='0'; e12 <='1'; e13 <='0'; e14 <='0'; e15 <='0'; e16 <='1'; e1 <='1'; e2 <='0'; wait for period;
            e11 <='1'; e12 <='1'; e13 <='0'; e14 <='0'; e15 <='0'; e16 <='1'; e1 <='1'; e2 <='0'; wait for period;
            e11 <='0'; e12 <='0'; e13 <='1'; e14 <='0'; e15 <='0'; e16 <='1'; e1 <='1'; e2 <='0'; wait for period;
            e11 <='1'; e12 <='0'; e13 <='1'; e14 <='0'; e15 <='0'; e16 <='1'; e1 <='1'; e2 <='0'; wait for period;
            e11 <='0'; e12 <='1'; e13 <='1'; e14 <='0'; e15 <='0'; e16 <='1'; e1 <='1'; e2 <='0'; wait for period;
            e11 <='1'; e12 <='1'; e13 <='1'; e14 <='0'; e15 <='0'; e16 <='1'; e1 <='1'; e2 <='0'; wait for period;
            e11 <='0'; e12 <='0'; e13 <='0'; e14 <='1'; e15 <='0'; e16 <='1'; e1 <='1'; e2 <='0'; wait for period;
            e11 <='1'; e12 <='0'; e13 <='0'; e14 <='1'; e15 <='0'; e16 <='1'; e1 <='1'; e2 <='0'; wait for period;
            e11 <='0'; e12 <='1'; e13 <='0'; e14 <='1'; e15 <='0'; e16 <='1'; e1 <='1'; e2 <='0'; wait for period;
            e11 <='1'; e12 <='1'; e13 <='0'; e14 <='1'; e15 <='0'; e16 <='1'; e1 <='1'; e2 <='0'; wait for period;
            e11 <='0'; e12 <='0'; e13 <='1'; e14 <='1'; e15 <='0'; e16 <='1'; e1 <='1'; e2 <='0'; wait for period;
            e11 <='1'; e12 <='0'; e13 <='1'; e14 <='1'; e15 <='0'; e16 <='1'; e1 <='1'; e2 <='0'; wait for period;
            e11 <='0'; e12 <='1'; e13 <='1'; e14 <='1'; e15 <='0'; e16 <='1'; e1 <='1'; e2 <='0'; wait for period;
            e11 <='1'; e12 <='1'; e13 <='1'; e14 <='1'; e15 <='0'; e16 <='1'; e1 <='1'; e2 <='0'; wait for period;
            e11 <='0'; e12 <='0'; e13 <='0'; e14 <='0'; e15 <='1'; e16 <='1'; e1 <='1'; e2 <='0'; wait for period;
            e11 <='1'; e12 <='0'; e13 <='0'; e14 <='0'; e15 <='1'; e16 <='1'; e1 <='1'; e2 <='0'; wait for period;
            e11 <='0'; e12 <='1'; e13 <='0'; e14 <='0'; e15 <='1'; e16 <='1'; e1 <='1'; e2 <='0'; wait for period;
            e11 <='1'; e12 <='1'; e13 <='0'; e14 <='0'; e15 <='1'; e16 <='1'; e1 <='1'; e2 <='0'; wait for period;
            e11 <='0'; e12 <='0'; e13 <='1'; e14 <='0'; e15 <='1'; e16 <='1'; e1 <='1'; e2 <='0'; wait for period;
            e11 <='1'; e12 <='0'; e13 <='1'; e14 <='0'; e15 <='1'; e16 <='1'; e1 <='1'; e2 <='0'; wait for period;
            e11 <='0'; e12 <='1'; e13 <='1'; e14 <='0'; e15 <='1'; e16 <='1'; e1 <='1'; e2 <='0'; wait for period;
            e11 <='1'; e12 <='1'; e13 <='1'; e14 <='0'; e15 <='1'; e16 <='1'; e1 <='1'; e2 <='0'; wait for period;
            e11 <='0'; e12 <='0'; e13 <='0'; e14 <='1'; e15 <='1'; e16 <='1'; e1 <='1'; e2 <='0'; wait for period;
            e11 <='1'; e12 <='0'; e13 <='0'; e14 <='1'; e15 <='1'; e16 <='1'; e1 <='1'; e2 <='0'; wait for period;
            e11 <='0'; e12 <='1'; e13 <='0'; e14 <='1'; e15 <='1'; e16 <='1'; e1 <='1'; e2 <='0'; wait for period;
            e11 <='1'; e12 <='1'; e13 <='0'; e14 <='1'; e15 <='1'; e16 <='1'; e1 <='1'; e2 <='0'; wait for period;
            e11 <='0'; e12 <='0'; e13 <='1'; e14 <='1'; e15 <='1'; e16 <='1'; e1 <='1'; e2 <='0'; wait for period;
            e11 <='1'; e12 <='0'; e13 <='1'; e14 <='1'; e15 <='1'; e16 <='1'; e1 <='1'; e2 <='0'; wait for period;
            e11 <='0'; e12 <='1'; e13 <='1'; e14 <='1'; e15 <='1'; e16 <='1'; e1 <='1'; e2 <='0'; wait for period;
            e11 <='1'; e12 <='1'; e13 <='1'; e14 <='1'; e15 <='1'; e16 <='1'; e1 <='1'; e2 <='0'; wait for period; -----
            e11 <='0'; e12 <='0'; e13 <='0'; e14 <='0'; e15 <='0'; e16 <='0'; e1 <='0'; e2 <='1'; wait for period;
            e11 <='1'; e12 <='0'; e13 <='0'; e14 <='0'; e15 <='0'; e16 <='0'; e1 <='0'; e2 <='1'; wait for period;
            e11 <='0'; e12 <='1'; e13 <='0'; e14 <='0'; e15 <='0'; e16 <='0'; e1 <='0'; e2 <='1'; wait for period;
            e11 <='1'; e12 <='1'; e13 <='0'; e14 <='0'; e15 <='0'; e16 <='0'; e1 <='0'; e2 <='1'; wait for period;
            e11 <='0'; e12 <='0'; e13 <='1'; e14 <='0'; e15 <='0'; e16 <='0'; e1 <='0'; e2 <='1'; wait for period;
            e11 <='1'; e12 <='0'; e13 <='1'; e14 <='0'; e15 <='0'; e16 <='0'; e1 <='0'; e2 <='1'; wait for period;
            e11 <='0'; e12 <='1'; e13 <='1'; e14 <='0'; e15 <='0'; e16 <='0'; e1 <='0'; e2 <='1'; wait for period;
            e11 <='1'; e12 <='1'; e13 <='1'; e14 <='0'; e15 <='0'; e16 <='0'; e1 <='0'; e2 <='1'; wait for period;
            e11 <='0'; e12 <='0'; e13 <='0'; e14 <='1'; e15 <='0'; e16 <='0'; e1 <='0'; e2 <='1'; wait for period;
            e11 <='1'; e12 <='0'; e13 <='0'; e14 <='1'; e15 <='0'; e16 <='0'; e1 <='0'; e2 <='1'; wait for period;
            e11 <='0'; e12 <='1'; e13 <='0'; e14 <='1'; e15 <='0'; e16 <='0'; e1 <='0'; e2 <='1'; wait for period;
            e11 <='1'; e12 <='1'; e13 <='0'; e14 <='1'; e15 <='0'; e16 <='0'; e1 <='0'; e2 <='1'; wait for period;
            e11 <='0'; e12 <='0'; e13 <='1'; e14 <='1'; e15 <='0'; e16 <='0'; e1 <='0'; e2 <='1'; wait for period;
            e11 <='1'; e12 <='0'; e13 <='1'; e14 <='1'; e15 <='0'; e16 <='0'; e1 <='0'; e2 <='1'; wait for period;
            e11 <='0'; e12 <='1'; e13 <='1'; e14 <='1'; e15 <='0'; e16 <='0'; e1 <='0'; e2 <='1'; wait for period;
            e11 <='1'; e12 <='1'; e13 <='1'; e14 <='1'; e15 <='0'; e16 <='0'; e1 <='0'; e2 <='1'; wait for period;
            e11 <='0'; e12 <='0'; e13 <='0'; e14 <='0'; e15 <='1'; e16 <='0'; e1 <='0'; e2 <='1'; wait for period;
            e11 <='1'; e12 <='0'; e13 <='0'; e14 <='0'; e15 <='1'; e16 <='0'; e1 <='0'; e2 <='1'; wait for period;
            e11 <='0'; e12 <='1'; e13 <='0'; e14 <='0'; e15 <='1'; e16 <='0'; e1 <='0'; e2 <='1'; wait for period;
            e11 <='1'; e12 <='1'; e13 <='0'; e14 <='0'; e15 <='1'; e16 <='0'; e1 <='0'; e2 <='1'; wait for period;
            e11 <='0'; e12 <='0'; e13 <='1'; e14 <='0'; e15 <='1'; e16 <='0'; e1 <='0'; e2 <='1'; wait for period;
            e11 <='1'; e12 <='0'; e13 <='1'; e14 <='0'; e15 <='1'; e16 <='0'; e1 <='0'; e2 <='1'; wait for period;
            e11 <='0'; e12 <='1'; e13 <='1'; e14 <='0'; e15 <='1'; e16 <='0'; e1 <='0'; e2 <='1'; wait for period;
            e11 <='1'; e12 <='1'; e13 <='1'; e14 <='0'; e15 <='1'; e16 <='0'; e1 <='0'; e2 <='1'; wait for period;
            e11 <='0'; e12 <='0'; e13 <='0'; e14 <='1'; e15 <='1'; e16 <='0'; e1 <='0'; e2 <='1'; wait for period;
            e11 <='1'; e12 <='0'; e13 <='0'; e14 <='1'; e15 <='1'; e16 <='0'; e1 <='0'; e2 <='1'; wait for period;
            e11 <='0'; e12 <='1'; e13 <='0'; e14 <='1'; e15 <='1'; e16 <='0'; e1 <='0'; e2 <='1'; wait for period;
            e11 <='1'; e12 <='1'; e13 <='0'; e14 <='1'; e15 <='1'; e16 <='0'; e1 <='0'; e2 <='1'; wait for period;
            e11 <='0'; e12 <='0'; e13 <='1'; e14 <='1'; e15 <='1'; e16 <='0'; e1 <='0'; e2 <='1'; wait for period;
            e11 <='1'; e12 <='0'; e13 <='1'; e14 <='1'; e15 <='1'; e16 <='0'; e1 <='0'; e2 <='1'; wait for period;
            e11 <='0'; e12 <='1'; e13 <='1'; e14 <='1'; e15 <='1'; e16 <='0'; e1 <='0'; e2 <='1'; wait for period;
            e11 <='1'; e12 <='1'; e13 <='1'; e14 <='1'; e15 <='1'; e16 <='0'; e1 <='0'; e2 <='1'; wait for period;
            e11 <='0'; e12 <='0'; e13 <='0'; e14 <='0'; e15 <='0'; e16 <='1'; e1 <='0'; e2 <='1'; wait for period;
            e11 <='1'; e12 <='0'; e13 <='0'; e14 <='0'; e15 <='0'; e16 <='1'; e1 <='0'; e2 <='1'; wait for period;
            e11 <='0'; e12 <='1'; e13 <='0'; e14 <='0'; e15 <='0'; e16 <='1'; e1 <='0'; e2 <='1'; wait for period;
            e11 <='1'; e12 <='1'; e13 <='0'; e14 <='0'; e15 <='0'; e16 <='1'; e1 <='0'; e2 <='1'; wait for period;
            e11 <='0'; e12 <='0'; e13 <='1'; e14 <='0'; e15 <='0'; e16 <='1'; e1 <='0'; e2 <='1'; wait for period;
            e11 <='1'; e12 <='0'; e13 <='1'; e14 <='0'; e15 <='0'; e16 <='1'; e1 <='0'; e2 <='1'; wait for period;
            e11 <='0'; e12 <='1'; e13 <='1'; e14 <='0'; e15 <='0'; e16 <='1'; e1 <='0'; e2 <='1'; wait for period;
            e11 <='1'; e12 <='1'; e13 <='1'; e14 <='0'; e15 <='0'; e16 <='1'; e1 <='0'; e2 <='1'; wait for period;
            e11 <='0'; e12 <='0'; e13 <='0'; e14 <='1'; e15 <='0'; e16 <='1'; e1 <='0'; e2 <='1'; wait for period;
            e11 <='1'; e12 <='0'; e13 <='0'; e14 <='1'; e15 <='0'; e16 <='1'; e1 <='0'; e2 <='1'; wait for period;
            e11 <='0'; e12 <='1'; e13 <='0'; e14 <='1'; e15 <='0'; e16 <='1'; e1 <='0'; e2 <='1'; wait for period;
            e11 <='1'; e12 <='1'; e13 <='0'; e14 <='1'; e15 <='0'; e16 <='1'; e1 <='0'; e2 <='1'; wait for period;
            e11 <='0'; e12 <='0'; e13 <='1'; e14 <='1'; e15 <='0'; e16 <='1'; e1 <='0'; e2 <='1'; wait for period;
            e11 <='1'; e12 <='0'; e13 <='1'; e14 <='1'; e15 <='0'; e16 <='1'; e1 <='0'; e2 <='1'; wait for period;
            e11 <='0'; e12 <='1'; e13 <='1'; e14 <='1'; e15 <='0'; e16 <='1'; e1 <='0'; e2 <='1'; wait for period;
            e11 <='1'; e12 <='1'; e13 <='1'; e14 <='1'; e15 <='0'; e16 <='1'; e1 <='0'; e2 <='1'; wait for period;
            e11 <='0'; e12 <='0'; e13 <='0'; e14 <='0'; e15 <='1'; e16 <='1'; e1 <='0'; e2 <='1'; wait for period;
            e11 <='1'; e12 <='0'; e13 <='0'; e14 <='0'; e15 <='1'; e16 <='1'; e1 <='0'; e2 <='1'; wait for period;
            e11 <='0'; e12 <='1'; e13 <='0'; e14 <='0'; e15 <='1'; e16 <='1'; e1 <='0'; e2 <='1'; wait for period;
            e11 <='1'; e12 <='1'; e13 <='0'; e14 <='0'; e15 <='1'; e16 <='1'; e1 <='0'; e2 <='1'; wait for period;
            e11 <='0'; e12 <='0'; e13 <='1'; e14 <='0'; e15 <='1'; e16 <='1'; e1 <='0'; e2 <='1'; wait for period;
            e11 <='1'; e12 <='0'; e13 <='1'; e14 <='0'; e15 <='1'; e16 <='1'; e1 <='0'; e2 <='1'; wait for period;
            e11 <='0'; e12 <='1'; e13 <='1'; e14 <='0'; e15 <='1'; e16 <='1'; e1 <='0'; e2 <='1'; wait for period;
            e11 <='1'; e12 <='1'; e13 <='1'; e14 <='0'; e15 <='1'; e16 <='1'; e1 <='0'; e2 <='1'; wait for period;
            e11 <='0'; e12 <='0'; e13 <='0'; e14 <='1'; e15 <='1'; e16 <='1'; e1 <='0'; e2 <='1'; wait for period;
            e11 <='1'; e12 <='0'; e13 <='0'; e14 <='1'; e15 <='1'; e16 <='1'; e1 <='0'; e2 <='1'; wait for period;
            e11 <='0'; e12 <='1'; e13 <='0'; e14 <='1'; e15 <='1'; e16 <='1'; e1 <='0'; e2 <='1'; wait for period;
            e11 <='1'; e12 <='1'; e13 <='0'; e14 <='1'; e15 <='1'; e16 <='1'; e1 <='0'; e2 <='1'; wait for period;
            e11 <='0'; e12 <='0'; e13 <='1'; e14 <='1'; e15 <='1'; e16 <='1'; e1 <='0'; e2 <='1'; wait for period;
            e11 <='1'; e12 <='0'; e13 <='1'; e14 <='1'; e15 <='1'; e16 <='1'; e1 <='0'; e2 <='1'; wait for period;
            e11 <='0'; e12 <='1'; e13 <='1'; e14 <='1'; e15 <='1'; e16 <='1'; e1 <='0'; e2 <='1'; wait for period;
            e11 <='1'; e12 <='1'; e13 <='1'; e14 <='1'; e15 <='1'; e16 <='1'; e1 <='0'; e2 <='1'; wait for period;
            e11 <='0'; e12 <='0'; e13 <='0'; e14 <='0'; e15 <='0'; e16 <='0'; e1 <='1'; e2 <='1'; wait for period;
            e11 <='1'; e12 <='0'; e13 <='0'; e14 <='0'; e15 <='0'; e16 <='0'; e1 <='1'; e2 <='1'; wait for period;
            e11 <='0'; e12 <='1'; e13 <='0'; e14 <='0'; e15 <='0'; e16 <='0'; e1 <='1'; e2 <='1'; wait for period;
            e11 <='1'; e12 <='1'; e13 <='0'; e14 <='0'; e15 <='0'; e16 <='0'; e1 <='1'; e2 <='1'; wait for period;
            e11 <='0'; e12 <='0'; e13 <='1'; e14 <='0'; e15 <='0'; e16 <='0'; e1 <='1'; e2 <='1'; wait for period;
            e11 <='1'; e12 <='0'; e13 <='1'; e14 <='0'; e15 <='0'; e16 <='0'; e1 <='1'; e2 <='1'; wait for period;
            e11 <='0'; e12 <='1'; e13 <='1'; e14 <='0'; e15 <='0'; e16 <='0'; e1 <='1'; e2 <='1'; wait for period;
            e11 <='1'; e12 <='1'; e13 <='1'; e14 <='0'; e15 <='0'; e16 <='0'; e1 <='1'; e2 <='1'; wait for period;
            e11 <='0'; e12 <='0'; e13 <='0'; e14 <='1'; e15 <='0'; e16 <='0'; e1 <='1'; e2 <='1'; wait for period;
            e11 <='1'; e12 <='0'; e13 <='0'; e14 <='1'; e15 <='0'; e16 <='0'; e1 <='1'; e2 <='1'; wait for period;
            e11 <='0'; e12 <='1'; e13 <='0'; e14 <='1'; e15 <='0'; e16 <='0'; e1 <='1'; e2 <='1'; wait for period;
            e11 <='1'; e12 <='1'; e13 <='0'; e14 <='1'; e15 <='0'; e16 <='0'; e1 <='1'; e2 <='1'; wait for period;
            e11 <='0'; e12 <='0'; e13 <='1'; e14 <='1'; e15 <='0'; e16 <='0'; e1 <='1'; e2 <='1'; wait for period;
            e11 <='1'; e12 <='0'; e13 <='1'; e14 <='1'; e15 <='0'; e16 <='0'; e1 <='1'; e2 <='1'; wait for period;
            e11 <='0'; e12 <='1'; e13 <='1'; e14 <='1'; e15 <='0'; e16 <='0'; e1 <='1'; e2 <='1'; wait for period;
            e11 <='1'; e12 <='1'; e13 <='1'; e14 <='1'; e15 <='0'; e16 <='0'; e1 <='1'; e2 <='1'; wait for period;
            e11 <='0'; e12 <='0'; e13 <='0'; e14 <='0'; e15 <='1'; e16 <='0'; e1 <='1'; e2 <='1'; wait for period;
            e11 <='1'; e12 <='0'; e13 <='0'; e14 <='0'; e15 <='1'; e16 <='0'; e1 <='1'; e2 <='1'; wait for period;
            e11 <='0'; e12 <='1'; e13 <='0'; e14 <='0'; e15 <='1'; e16 <='0'; e1 <='1'; e2 <='1'; wait for period;
            e11 <='1'; e12 <='1'; e13 <='0'; e14 <='0'; e15 <='1'; e16 <='0'; e1 <='1'; e2 <='1'; wait for period;
            e11 <='0'; e12 <='0'; e13 <='1'; e14 <='0'; e15 <='1'; e16 <='0'; e1 <='1'; e2 <='1'; wait for period;
            e11 <='1'; e12 <='0'; e13 <='1'; e14 <='0'; e15 <='1'; e16 <='0'; e1 <='1'; e2 <='1'; wait for period;
            e11 <='0'; e12 <='1'; e13 <='1'; e14 <='0'; e15 <='1'; e16 <='0'; e1 <='1'; e2 <='1'; wait for period;
            e11 <='1'; e12 <='1'; e13 <='1'; e14 <='0'; e15 <='1'; e16 <='0'; e1 <='1'; e2 <='1'; wait for period;
            e11 <='0'; e12 <='0'; e13 <='0'; e14 <='1'; e15 <='1'; e16 <='0'; e1 <='1'; e2 <='1'; wait for period;
            e11 <='1'; e12 <='0'; e13 <='0'; e14 <='1'; e15 <='1'; e16 <='0'; e1 <='1'; e2 <='1'; wait for period;
            e11 <='0'; e12 <='1'; e13 <='0'; e14 <='1'; e15 <='1'; e16 <='0'; e1 <='1'; e2 <='1'; wait for period;
            e11 <='1'; e12 <='1'; e13 <='0'; e14 <='1'; e15 <='1'; e16 <='0'; e1 <='1'; e2 <='1'; wait for period;
            e11 <='0'; e12 <='0'; e13 <='1'; e14 <='1'; e15 <='1'; e16 <='0'; e1 <='1'; e2 <='1'; wait for period;
            e11 <='1'; e12 <='0'; e13 <='1'; e14 <='1'; e15 <='1'; e16 <='0'; e1 <='1'; e2 <='1'; wait for period;
            e11 <='0'; e12 <='1'; e13 <='1'; e14 <='1'; e15 <='1'; e16 <='0'; e1 <='1'; e2 <='1'; wait for period;
            e11 <='1'; e12 <='1'; e13 <='1'; e14 <='1'; e15 <='1'; e16 <='0'; e1 <='1'; e2 <='1'; wait for period;
            e11 <='0'; e12 <='0'; e13 <='0'; e14 <='0'; e15 <='0'; e16 <='1'; e1 <='1'; e2 <='1'; wait for period;
            e11 <='1'; e12 <='0'; e13 <='0'; e14 <='0'; e15 <='0'; e16 <='1'; e1 <='1'; e2 <='1'; wait for period;
            e11 <='0'; e12 <='1'; e13 <='0'; e14 <='0'; e15 <='0'; e16 <='1'; e1 <='1'; e2 <='1'; wait for period;
            e11 <='1'; e12 <='1'; e13 <='0'; e14 <='0'; e15 <='0'; e16 <='1'; e1 <='1'; e2 <='1'; wait for period;
            e11 <='0'; e12 <='0'; e13 <='1'; e14 <='0'; e15 <='0'; e16 <='1'; e1 <='1'; e2 <='1'; wait for period;
            e11 <='1'; e12 <='0'; e13 <='1'; e14 <='0'; e15 <='0'; e16 <='1'; e1 <='1'; e2 <='1'; wait for period;
            e11 <='0'; e12 <='1'; e13 <='1'; e14 <='0'; e15 <='0'; e16 <='1'; e1 <='1'; e2 <='1'; wait for period;
            e11 <='1'; e12 <='1'; e13 <='1'; e14 <='0'; e15 <='0'; e16 <='1'; e1 <='1'; e2 <='1'; wait for period;
            e11 <='0'; e12 <='0'; e13 <='0'; e14 <='1'; e15 <='0'; e16 <='1'; e1 <='1'; e2 <='1'; wait for period;
            e11 <='1'; e12 <='0'; e13 <='0'; e14 <='1'; e15 <='0'; e16 <='1'; e1 <='1'; e2 <='1'; wait for period;
            e11 <='0'; e12 <='1'; e13 <='0'; e14 <='1'; e15 <='0'; e16 <='1'; e1 <='1'; e2 <='1'; wait for period;
            e11 <='1'; e12 <='1'; e13 <='0'; e14 <='1'; e15 <='0'; e16 <='1'; e1 <='1'; e2 <='1'; wait for period;
            e11 <='0'; e12 <='0'; e13 <='1'; e14 <='1'; e15 <='0'; e16 <='1'; e1 <='1'; e2 <='1'; wait for period;
            e11 <='1'; e12 <='0'; e13 <='1'; e14 <='1'; e15 <='0'; e16 <='1'; e1 <='1'; e2 <='1'; wait for period;
            e11 <='0'; e12 <='1'; e13 <='1'; e14 <='1'; e15 <='0'; e16 <='1'; e1 <='1'; e2 <='1'; wait for period;
            e11 <='1'; e12 <='1'; e13 <='1'; e14 <='1'; e15 <='0'; e16 <='1'; e1 <='1'; e2 <='1'; wait for period;
            e11 <='0'; e12 <='0'; e13 <='0'; e14 <='0'; e15 <='1'; e16 <='1'; e1 <='1'; e2 <='1'; wait for period;
            e11 <='1'; e12 <='0'; e13 <='0'; e14 <='0'; e15 <='1'; e16 <='1'; e1 <='1'; e2 <='1'; wait for period;
            e11 <='0'; e12 <='1'; e13 <='0'; e14 <='0'; e15 <='1'; e16 <='1'; e1 <='1'; e2 <='1'; wait for period;
            e11 <='1'; e12 <='1'; e13 <='0'; e14 <='0'; e15 <='1'; e16 <='1'; e1 <='1'; e2 <='1'; wait for period;
            e11 <='0'; e12 <='0'; e13 <='1'; e14 <='0'; e15 <='1'; e16 <='1'; e1 <='1'; e2 <='1'; wait for period;
            e11 <='1'; e12 <='0'; e13 <='1'; e14 <='0'; e15 <='1'; e16 <='1'; e1 <='1'; e2 <='1'; wait for period;
            e11 <='0'; e12 <='1'; e13 <='1'; e14 <='0'; e15 <='1'; e16 <='1'; e1 <='1'; e2 <='1'; wait for period;
            e11 <='1'; e12 <='1'; e13 <='1'; e14 <='0'; e15 <='1'; e16 <='1'; e1 <='1'; e2 <='1'; wait for period;
            e11 <='0'; e12 <='0'; e13 <='0'; e14 <='1'; e15 <='1'; e16 <='1'; e1 <='1'; e2 <='1'; wait for period;
            e11 <='1'; e12 <='0'; e13 <='0'; e14 <='1'; e15 <='1'; e16 <='1'; e1 <='1'; e2 <='1'; wait for period;
            e11 <='0'; e12 <='1'; e13 <='0'; e14 <='1'; e15 <='1'; e16 <='1'; e1 <='1'; e2 <='1'; wait for period;
            e11 <='1'; e12 <='1'; e13 <='0'; e14 <='1'; e15 <='1'; e16 <='1'; e1 <='1'; e2 <='1'; wait for period;
            e11 <='0'; e12 <='0'; e13 <='1'; e14 <='1'; e15 <='1'; e16 <='1'; e1 <='1'; e2 <='1'; wait for period;
            e11 <='1'; e12 <='0'; e13 <='1'; e14 <='1'; e15 <='1'; e16 <='1'; e1 <='1'; e2 <='1'; wait for period;
            e11 <='0'; e12 <='1'; e13 <='1'; e14 <='1'; e15 <='1'; e16 <='1'; e1 <='1'; e2 <='1'; wait for period;
            e11 <='1'; e12 <='1'; e13 <='1'; e14 <='1'; e15 <='1'; e16 <='1'; e1 <='1'; e2 <='1'; wait for period;
            e11 <='0'; e12 <='0'; e13 <='0'; e14 <='0'; e15 <='0'; e16 <='0'; e1 <='0'; e2 <='0'; wait;
        end process;
        
    Transmit : Main PORT MAP(e1, e2, e11, e12, e13, e14, e15, e16, l1, l2, l11, l12, l13, l14, l15, l16, a, b, c, d, e, f, g, dp);
end Behavioral;
