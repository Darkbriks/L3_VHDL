library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity Gate_Nand is
    Port ( e1 : in STD_LOGIC;
           e2 : in STD_LOGIC;
           res : out std_logic);
end Gate_Nand;

architecture Behavioral of Gate_Nand is

begin
    res<='1' when not (e1='1' and e2='1') else '0';
end Behavioral;
